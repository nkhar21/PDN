*

.SUBCKT		b4_1_092725_171600_21104
+			decap_port1_1
+			decap_port1_2
+			decap_port2_1
+			decap_port2_2
+			ic_port_1
+			ic_port_2
*The following is the Cadence MCP(model connection protocol) Section
***********************************
*[MCP Begin]
*[MCP Ver] 1.1
*[MCP Source] Cadence Design Systems, Inc. Layout Workbench 24.1.0.10141.541387   000 9/27/2025
*
***********************************
*
*[REM]The following is the info for component connection decap_port1
*[REM]**********************************
*[Connection] decap_port1 cap 2
*[Power Nets]
*1	decap_port1_1	pwr	0.0250000	0.0300000
*[Ground Nets]
*2	decap_port1_2	gnd	0.0280000	0.0300000
*[Signal Nets]
*
*[REM]The following is the info for component connection decap_port2
*[REM]**********************************
*[Connection] decap_port2 cap 2
*[Power Nets]
*1	decap_port2_1	pwr	0.0250000	0.0250000
*[Ground Nets]
*2	decap_port2_2	gnd	0.0280000	0.0250000
*[Signal Nets]
*
*[REM]The following is the info for component connection ic_port
*[REM]**********************************
*[Connection] ic_port ic 2
*[Power Nets]
*1	ic_port_1	pwr	0.0350000	0.0350000
*[Ground Nets]
*2	ic_port_2	gnd	0.0350000	0.0300000
*[Signal Nets]
*
*[MCP End]
*
*This concludes the MCP section
*Define the S element, the Model file is output from BNP

.MODEL   Spara   S		
+		BNPFILE = "b4_1_092725_171600_21104.bnp"

S		
+			decap_port1_1	decap_port1_2
+			decap_port2_1	decap_port2_2
+			ic_port_1	ic_port_2
+			MNAME = Spara

*
.ENDS
*
*
